library verilog;
use verilog.vl_types.all;
entity p4_tb1 is
end p4_tb1;
