library verilog;
use verilog.vl_types.all;
entity circuit_02 is
    port(
        y2              : out    vl_logic;
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        x4              : in     vl_logic
    );
end circuit_02;
