library verilog;
use verilog.vl_types.all;
entity circuit_01 is
    port(
        y               : out    vl_logic;
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic
    );
end circuit_01;
