library verilog;
use verilog.vl_types.all;
entity circuit_tb1 is
end circuit_tb1;
