library verilog;
use verilog.vl_types.all;
entity circuit_01_tb1 is
end circuit_01_tb1;
